module lab6(input logic inLED,
            ouput logic outLED);
    assign outLED = inLED;
endmodule